library verilog;
use verilog.vl_types.all;
entity tb is
    generic(
        n               : integer := 9
    );
end tb;
