library verilog;
use verilog.vl_types.all;
entity tb is
    generic(
        N               : integer := 4
    );
end tb;
