module modulus_operator(x,y,out);
input [3:0] x,y;
output [3:0] out;
	assign out=x%y;
endmodule
	
