library verilog;
use verilog.vl_types.all;
entity tb is
    generic(
        S               : integer := 2;
        M               : integer := 3
    );
end tb;
