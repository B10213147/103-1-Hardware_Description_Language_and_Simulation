library verilog;
use verilog.vl_types.all;
entity tb is
    generic(
        N               : integer := 5
    );
end tb;
